
//* ----- Global parameters -----
`define HAP_MAX_LENGTH              128
`define READ_MAX_LENGTH             64

//* DP for Genotyping
`define DP_PAIRHMM_SCORE_BITWIDTH   16

`define CONST_M2M                   -1
`define CONST_M2I                   -3072
`define CONST_I2I                   -1024
`define CONST_I2M                   -47

`define CONST_MATCH_BITWIDTH        16
`define CONST_BQ0_MATCH_SCORE       -443
`define CONST_BQ1_MATCH_SCORE       -37
`define CONST_BQ2_MATCH_SCORE       -1
`define CONST_BQ3_MATCH_SCORE       0

`define CONST_MISMATCH_BITWIDTH     16
`define CONST_BQ0_MISMATCH_SCORE    -4276
`define CONST_BQ1_MISMATCH_SCORE    -3043
`define CONST_BQ2_MISMATCH_SCORE    -1615
`define CONST_BQ3_MISMATCH_SCORE    -693



`define AVALON_RS232_BASE_ADDR  5'h00

